** sch_path: /workspaces/Talleres-fork/resuelto-klayout/schematic/inv.sch

.subckt inv vout vdd vin vss
*.PININFO vout:B vdd:B vin:B vss:B
XM1 vout vin vdd vdd pfet_03v3 L=0.280u W=0.720u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 vout vin vss vss nfet_03v3 L=0.280u W=0.360u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends
.end
