*************************************************
* Tools: LTspice + L-Edit(layout)				*
*************************************************

* Models
.include "2um_CMOS.modlib"

* Dise�o de inversor unitario con informacion de layout
.subckt unit_inv In Out1 Vdd Vss
* Transistores CMOS
* MOSFET Syntax: Mxxx Nd Ng Ns Nb <model>
M5 Vdd In Out1 Vdd P_2u L=2u W=6u AD=72p PD=48u AS=36p PS=24u
M6 Out1 In Vdd Vdd P_2u L=2u W=6u AD=36p PD=24u AS=72p PS=48u
M7 Out1 In Vss Vss N_2u L=2u W=6u AD=36p PD=24u AS=36p PS=24u
* Capacitancias parasitas
Cpar1 Vdd 0 441.28174f
Cpar2 Vss 0 310.12743f
Cpar3 In 0 10.420182f
Cpar4 Out1 0 139.14517f
.ends

******************
* Retardo de propagacion inversor unitario
* Voltage sources
V_dd V_dd 0 DC 5
* Vxxx n+ n- PULSE(V1 V2 Tdelay Trise Tfall Ton Tperiod Ncycles
V_in V_in 0 PULSE(0 5 1n 0p1 0p1 5n 10n)
* Instancias de sub-circuitos
X V_in Vout V_dd 0 unit_inv
* Capacitancias de carga
CL Vout_unit 0 83.361456f
* Analysis
.tran 12n


.backanno
.end
