magic
tech sky130A
timestamp 1685238938
<< nwell >>
rect 0 250 280 500
<< nmos >>
rect 125 60 155 210
<< pmos >>
rect 55 270 85 420
rect 125 270 155 420
rect 195 270 225 420
<< ndiff >>
rect 90 195 125 210
rect 90 75 95 195
rect 115 75 125 195
rect 90 60 125 75
rect 155 195 190 210
rect 155 75 165 195
rect 185 75 190 195
rect 155 60 190 75
<< pdiff >>
rect 20 405 55 420
rect 20 285 25 405
rect 45 285 55 405
rect 20 270 55 285
rect 85 405 125 420
rect 85 285 95 405
rect 115 285 125 405
rect 85 270 125 285
rect 155 405 195 420
rect 155 285 165 405
rect 185 285 195 405
rect 155 270 195 285
rect 225 405 260 420
rect 225 285 235 405
rect 255 285 260 405
rect 225 270 260 285
<< ndiffc >>
rect 95 75 115 195
rect 165 75 185 195
<< pdiffc >>
rect 25 285 45 405
rect 95 285 115 405
rect 165 285 185 405
rect 235 285 255 405
<< psubdiff >>
rect 20 25 260 30
rect 20 5 35 25
rect 245 5 260 25
rect 20 0 260 5
<< nsubdiff >>
rect 20 475 260 480
rect 20 455 35 475
rect 245 455 260 475
rect 20 450 260 455
<< psubdiffcont >>
rect 35 5 245 25
<< nsubdiffcont >>
rect 35 455 245 475
<< poly >>
rect 55 420 85 435
rect 125 420 155 435
rect 195 420 225 435
rect 55 255 85 270
rect 30 250 85 255
rect 125 250 155 270
rect 195 250 225 270
rect 30 245 225 250
rect 30 225 40 245
rect 60 225 225 245
rect 30 220 225 225
rect 30 215 70 220
rect 125 210 155 220
rect 125 45 155 60
<< polycont >>
rect 40 225 60 245
<< locali >>
rect 0 475 280 480
rect 0 455 35 475
rect 245 455 280 475
rect 0 450 280 455
rect 25 415 45 450
rect 165 415 185 450
rect 20 405 50 415
rect 20 285 25 405
rect 45 285 50 405
rect 20 275 50 285
rect 90 405 120 415
rect 90 285 95 405
rect 115 285 120 405
rect 90 275 120 285
rect 160 405 190 415
rect 160 285 165 405
rect 185 285 190 405
rect 160 275 190 285
rect 230 405 260 415
rect 230 285 235 405
rect 255 285 260 405
rect 230 275 260 285
rect 30 245 70 255
rect 0 225 40 245
rect 60 225 70 245
rect 95 245 115 275
rect 235 245 255 275
rect 95 225 280 245
rect 30 215 70 225
rect 165 205 185 225
rect 90 195 120 205
rect 90 75 95 195
rect 115 75 120 195
rect 90 65 120 75
rect 160 195 190 205
rect 160 75 165 195
rect 185 75 190 195
rect 160 65 190 75
rect 95 30 115 65
rect 0 25 280 30
rect 0 5 35 25
rect 245 5 280 25
rect 0 0 280 5
<< labels >>
rlabel locali 260 225 280 245 3 Vout
rlabel locali 0 225 20 245 7 Vin
rlabel locali 0 5 20 25 5 Gnd
rlabel locali 0 455 20 475 1 Vdd
<< end >>
