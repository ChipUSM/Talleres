* Extracted by KLayout with SG13G2 LVS runset on : 19/05/2025 19:27

.SUBCKT inv Vin Vdd Vss Vout
M$1 Vdd Vin Vout Vdd sg13_lv_pmos L=0.13u W=0.81u AS=0.2754p AD=0.2754p PS=2.3u
+ PD=2.3u
M$2 Vss Vin Vout Vss sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u
+ PD=1.28u
.ENDS inv
