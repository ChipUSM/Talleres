* NGSPICE file created from inv_flat.ext - technology: sky130A

.subckt inv_flat
X0 Vdd Vin Vout Vdd sky130_fd_pr__pfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.3
X1 Vout Vin Gnd Gnd sky130_fd_pr__nfet_01v8 ad=0.525 pd=3.7 as=0.525 ps=3.7 w=1.5 l=0.3
X2 Vout Vin Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0.3 pd=1.9 as=0.525 ps=3.7 w=1.5 l=0.3
X3 Vout Vin Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0.525 pd=3.7 as=0.3 ps=1.9 w=1.5 l=0.3
C0 Vdd Vout 0.306583f
C1 Vin Vdd 0.331762f
C2 Vin Vout 0.224963f
C3 Vout Gnd 0.301175f
C4 Vin Gnd 0.512965f
C5 Vdd Gnd 0.978789f
.ends

