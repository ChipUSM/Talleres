*

.include "2um_CMOS.modlib"
* MOSFET Syntax: Mxxx Nd Ng Ns Nb <model>

* NMOS with parasitic capacitances
.subckt nmos_parasitics D G S
M1 D G S S N_2u L=2u W=20u AD=110p PD=51u AS=110p PS=51u
Cpar1 S 0 333.96838f
Cpar2 G 0 6.824306f
Cpar3 D 0 208.80869f
.end

* NMOS 2 fingers, with parasitic capacitances
.subckt nmos_2fingers_parasitics D G S
M1 S G D S N_2u L=2u W=10u AD=110p PD=62u AS=60p PS=32u
M2 D G S S N_2u L=2u W=10u AD=60p PD=32u AS=110p PS=62u
Cpar1 S 0 410.68277f
Cpar2 D 0 114.3739f
Cpar3 G 0 8.2251705f
.end


* NMOS
R0 VDD D0 10k
M0 D0 G 0 0 N_2u L=2u W=20u
Cload0 D0 0 100f

R1 VDD D1 10k
X1 D1 G 0 nmos_parasitics
Cload1 D1 0 100f

R2 VDD D2 10k
X2 D2 G 0 nmos_2fingers_parasitics
Cload3 D2 GND 100f

Vdd VDD GND 5
* Vxx n+ n- PULSE(V1 V2 Tdelay Trise Tfall Ton Tperiod Ncycles
Vgs G GND PULSE(0 5 0.2n 1f 1f 10n 20n 1)
.tran 1n

.end
